Library IEEE;
use IEEE.std_logic_1164.all;
ENTITY sete_seg_bomba is
port(
	entrada_seg	:in std_logic_vector(5 downto 0);
	saida_seg :out std_logic_vector(0 to 13)
	);
end sete_seg_bomba;

ARCHITECTURE arc_seg of sete_seg_bomba is
begin
	with entrada_seg select
	saida_seg <="00000010000001" when "000000",		--0
				"00000011001111" when "000001",		--1
				"00000010010010" when "000010",		--2
				"00000010000110" when "000011",		--3
				"00000011001100" when "000100",		--4
				"00000010100100" when "000101",		--5
				"00000010100000" when "000110",		--6
				"00000010001111" when "000111",		--7
				"00000010000000" when "001000",		--8
				"00000010000100" when "001001",		--9
				"10011110000001" when "001010",		--10
				"10011111001111" when "001011",		--11
				"10011110010010" when "001100",		--12
				"10011110000110" when "001101",		--13
				"10011111001100" when "001110",		--14
				"10011110100100" when "001111",		--15
				"10011110100000" when "010000",		--16
				"10011110001111" when "010001",		--17
				"10011110000000" when "010010",		--18
				"10011110000100" when "010011",		--19
				"00100100000001" when "010100",		--20
				"00100101001111" when "010101",		--21
				"00100100010010" when "010110",		--22
				"00100100000110" when "010111",		--23
				"00100101001100" when "011000",		--24
				"00100100100100" when "011001",		--25
				"00100100100000" when "011010",		--26
				"00100100001111" when "011011",		--27
				"00100100000000" when "011100",		--28
				"00100100000100" when "011101",		--29
				"00001100000001" when "011110",		--30
				"00001101001111" when "011111",		--31
				"00001100010010" when "100000",		--32
				"00001100000110" when "100001",		--33
				"00001101001100" when "100010",		--34
				"00001100100100" when "100011",		--35
				"00001100100000" when "100100",		--36
				"00001100001111" when "100101",		--37
				"00001100000000" when "100110",		--38
				"00001100000100" when "100111",		--39
				"10011000000001" when "101000",		--40
				"10011001001111" when "101001",		--41
				"10011000010010" when "101010",		--42
				"10011000000110" when "101011",		--43
				"10011001001100" when "101100",		--44
				"10011000100100" when "101101",		--45
				"10011000100000" when "101110",		--46
				"10011000001111" when "101111",		--47
				"10011000000000" when "110000",		--48
				"10011000000100" when "110001",		--49
				"01001000000001" when "110010",		--50
				"01001001001111" when "110011",		--51
				"01001000010010" when "110100",		--52
				"01001000000110" when "110101",		--53
				"01001001001100" when "110110",		--54
				"01001000100100" when "110111",		--55
				"01001000100000" when "111000",		--56
				"01001000001111" when "111001",		--57
				"01001000000000" when "111010",		--58
				"01001000000100" when "111011",		--59
				"01000000000001" when "111100",		--60
				"01000000000001" when "111101",		--mantem o 60, quando 61
				"01000000000001" when "111110",		--mantem o 60, quando 62
				"01000000000001" when "111111",		--mantem o 60, quando 63
				"00000010000001" when others;
	
end arc_seg;
